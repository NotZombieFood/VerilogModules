module Excercise3(

	input [3:0] a,  //a son los switches 3-0
	input [3:0] b,  //b son los switches 15-11
	input ci,		 //cin es el switch 10
	output [6:0] display,
	output cout
);

wire co1,co2,co3;
wire [3:0] s;

FullAdder fa1 (
	.ci(ci),
	.a(a[0]),
	.b(b[0]),
	.s(s[0]),
	.co(co1)
);

FullAdder fa2 (
	.ci(co1),
	.a(a[1]),
	.b(b[1]),
	.s(s[1]),
	.co(co2)
);

FullAdder fa3 (
	.ci(co2),
	.a(a[2]),
	.b(b[2]),
	.s(s[2]),
	.co(co3)
);

FullAdder fa4 (
	.ci(co3),
	.a(a[3]),
	.b(b[3]),
	.s(s[3]),
	.co(cout)
);
/*
	assign display[0] = (s[3] & ~s[2] & ~s[1]) + (~s[3] & s[2] & s[0]) + (~s[3] & s[1]);
	assign display[1] = ( ~s[3] & s[2] & ~s[1] & ~s[0]) + ( s[3] & ~s[2] & ~s[1] ) + ( ~s[3] & ~s[2] & s[1] ) + ( ~s[3] & s[1] & s[0] );
	assign display[2] = (s[3] & ~s[2] & ~s[1] ) + (~s[3] & s[2] ) + (~s[3] & s[0] );
	assign display[3] = (s[3] & ~s[2] & ~s[1] & ~s[0] ) + (~s[3] & s[2] & ~s[1] & s[0] ) + ( ~s[3] & ~s[2] & s[1] ) + ( ~s[3] & s[1] & ~s[0] );
	assign display[4] = (s[3] & ~s[2] & ~s[1] & ~s[0] ) + ( ~s[3] & s[1] & ~s[0] );
	assign display[5] = (s[3] & ~s[2] & ~s[1] ) + ( ~s[3] & s[2] & ~s[1] ) + ( ~s[3] & s[2] & s[1] & ~s[0] );
	assign display[6] = (s[3] & ~s[2] & ~s[1] ) + ( ~s[3] & s[2] & ~s[1] ) + ( ~s[3] & ~s[2] & s[1] ) + ( ~s[2] & s[1] & ~s[0] );
*/




//													0											2										3												5
	assign display[0]= ((~s[3])&(~s[2])&(~s[1])&(~s[0]))|((~s[3])&(~s[2])&(s[1])&(~s[0]))|((~s[3])&(~s[2])&(s[1])&(s[0]))|((~s[3])&(s[2])&(~s[1])&(s[0]))|  ((~s[3])&(s[2])&(s[1])&(~s[0]))|((~s[3])&(s[2])&(s[1])&(s[0]))|((s[3])&(~s[2])&(~s[1])&(~s[0]))|((s[3])&(~s[2])&(~s[1])&(s[0]));
//					6											7										8											9			


//													0												1										2										3
	assign display[1]= ((~s[3])&(~s[2])&(~s[1])&(~s[0]))|((~s[3])&(~s[2])&(~s[1])&(s[0]))|((~s[3])&(~s[2])&(s[1])&(~s[0]))|((~s[3])&(~s[2])&(s[1])&(s[0]))| ((~s[3])&(s[2])&(~s[1])&(~s[0]))|((~s[3])&(s[2])&(s[1])&(s[0]))|((s[3])&(~s[2])&(~s[1])&(~s[0]))|((s[3])&(~s[2])&(~s[1])&(s[0]));	
//					4											7											8											9


//													0											1										3												4
	assign display[2]= ((~s[3])&(~s[2])&(~s[1])&(~s[0]))|((~s[3])&(~s[2])&(~s[1])&(s[0]))|((~s[3])&(~s[2])&(s[1])&(s[0]))|((~s[3])&(s[2])&(~s[1])&(~s[0]))|  ((~s[3])&(s[2])&(~s[1])&(s[0]))|((~s[3])&(s[2])&(s[1])&(~s[0]))|((~s[3])&(s[2])&(s[1])&(s[0]))|((s[3])&(~s[2])&(~s[1])&(~s[0]))|
//					5											6											7											8
	((s[3])&(~s[2])&(~s[1])&(s[0]));
//						9
	
	
//													0											2											3										5
	assign display[3]= ((~s[3])&(~s[2])&(~s[1])&(~s[0]))|((~s[3])&(~s[2])&(s[1])&(~s[0]))|((~s[3])&(~s[2])&(s[1])&(s[0]))|((~s[3])&(s[2])&(~s[1])&(s[0]))|  ((~s[3])&(s[2])&(s[1])&(~s[0]))|((s[3])&(~s[2])&(~s[1])&(~s[0]))|((s[3])&(~s[2])&(~s[1])&(s[0]));
//					6										8											9
	

//													0											2										6												8
	assign display[4]= ((~s[3])&(~s[2])&(~s[1])&(~s[0]))|((~s[3])&(~s[2])&(s[1])&(~s[0]))|((~s[3])&(s[2])&(s[1])&(~s[0]))|((s[3])&(~s[2])&(~s[1])&(~s[0]));


//													0												4										5							   			6
	assign display[5]= ((~s[3])&(~s[2])&(~s[1])&(~s[0]))|((~s[3])&(s[2])&(~s[1])&(~s[0]))|((~s[3])&(s[2])&(~s[1])&(s[0]))|(~(s[3])&(s[2])&(s[1])&(~s[0]))| ((s[3])&(~s[2])&(~s[1])&(~s[0]))|((s[3])&(~s[2])&(~s[1])&(s[0]));	
//					8											9


//													2										3												4										5
	assign display[6]= ((~s[3])&(~s[2])&(s[1])&(~s[0]))|((~s[3])&(~s[2])&(s[1])&(s[0]))|((~s[3])&(s[2])&(~s[1])&(~s[0]))|((~s[3])&(s[2])&(~s[1])&(s[0]))|((~s[3])&(s[2])&(s[1])&(~s[0]))|((s[3])&(~s[2])&(~s[1])&(~s[0]))|((s[3])&(~s[2])&(~s[1])&(s[0]));
//					6							8											9

	
endmodule